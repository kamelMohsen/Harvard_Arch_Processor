LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


