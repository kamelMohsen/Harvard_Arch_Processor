LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;



ENTITY BOB_EX_MEM IS
	PORT (
    RESET,STALL,CLK: IN STD_LOGIC;
    RESULT_IN, DESTINATION_IN,READ1_IN: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    WB_IN: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    MEM_IN: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
	FLAGS_IN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	INST_0_8_IN: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
	EFFECTIVE_ADDRESS_IN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	RESULT_OUT, DESTINATION_OUT,READ1_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    WB_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    MEM_OUT: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
	FLAGS_OUT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	INST_0_8_OUT: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
	EFFECTIVE_ADDRESS_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY BOB_EX_MEM;


ARCHITECTURE BOB_EX_MEM_ARCH OF BOB_EX_MEM IS
  

    --THE EX/MEM INST_0_8 Register  
    COMPONENT BOB_EX_MEM_INST_0_8 IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
	d : IN std_logic_vector(8 DOWNTO 0);
    q : OUT std_logic_vector(8 DOWNTO 0));
    
    END COMPONENT;

    --THE EX/MEM DESTINATION Register  
    COMPONENT BOB_EX_MEM_DESTINATION IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
	d : IN std_logic_vector(31 DOWNTO 0);
    q : OUT std_logic_vector(31 DOWNTO 0));
    
    END COMPONENT;

    --THE EX/MEM EFEECTIVE ADDRESS Register  
    COMPONENT BOB_EX_MEM_EFFECTIVE_ADDRESS IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
    d : IN std_logic_vector(15 DOWNTO 0);
    q : OUT std_logic_vector(15 DOWNTO 0));

    END COMPONENT;

    --THE EX/MEM WB Register  
    COMPONENT BOB_EX_MEM_WB IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
    d : IN std_logic_vector(4 DOWNTO 0);
    q : OUT std_logic_vector(4 DOWNTO 0));

    END COMPONENT;

    --THE EX/MEM MEM Register  
    COMPONENT BOB_EX_MEM_MEM IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
    d : IN std_logic_vector(8 DOWNTO 0);
    q : OUT std_logic_vector(8 DOWNTO 0));

    END COMPONENT;



    --THE EX/MEM RESULT Register  
    COMPONENT BOB_EX_MEM_RESULT IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
    d : IN std_logic_vector(31 DOWNTO 0);
    q : OUT std_logic_vector(31 DOWNTO 0));

    END COMPONENT;

    --THE EX/MEM FLAGS Register  
    COMPONENT BOB_EX_MEM_FLAGS IS 

    PORT(
    Clk,Rst,enable : IN std_logic;
    d : IN std_logic_vector(3 DOWNTO 0);
    q : OUT std_logic_vector(3 DOWNTO 0));

    END COMPONENT;



    SIGNAL NOT_STALL: STD_LOGIC;
    BEGIN	
    

    NOT_STALL <= NOT STALL;

	--THE WB Register
	EX_MEM_WB: BOB_EX_MEM_WB PORT MAP (CLK, RESET, NOT_STALL, WB_IN, WB_OUT);

	--THE MEM Register
	EX_MEM_MEM: BOB_EX_MEM_MEM PORT MAP (CLK, RESET, NOT_STALL, MEM_IN, MEM_OUT);

	--THE FALGS Register
	EX_MEM_FLAGS: BOB_EX_MEM_FLAGS PORT MAP (CLK, RESET, NOT_STALL, FLAGS_IN, FLAGS_OUT);

    --THE INST_0_8 Register
    EX_MEM_INST_0_8: BOB_EX_MEM_INST_0_8 PORT MAP (CLK, RESET, NOT_STALL, INST_0_8_IN, INST_0_8_OUT);

    --THE RESULT Register
    EX_MEM_RESULT: BOB_EX_MEM_RESULT PORT MAP (CLK, RESET, NOT_STALL, RESULT_IN, RESULT_OUT);

    --THE EFFECTIVE ADDRESS Register
	EX_MEM_EFFECTIVE_ADDRESS: BOB_EX_MEM_EFFECTIVE_ADDRESS PORT MAP (CLK, RESET, NOT_STALL, EFFECTIVE_ADDRESS_IN, EFFECTIVE_ADDRESS_OUT);
	
   --THE DESTINATION Register
    EX_MEM_DESTINATION: BOB_EX_MEM_DESTINATION PORT MAP (CLK, RESET, NOT_STALL, DESTINATION_IN, DESTINATION_OUT);

    --THE READ1 Register
    EX_MEM_READ1: BOB_EX_MEM_RESULT PORT MAP (CLK, RESET, NOT_STALL, READ1_IN, READ1_OUT);



    
END BOB_EX_MEM_ARCH;