LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ORR IS
 	PORT ( Input0, Input1 :IN STD_LOGIC; 
	Output0: OUT STD_LOGIC
	);
END ENTITY ORR;


ARCHITECTURE ORING OF ORR IS
BEGIN
	Output0 <= '1' WHEN Input0 ='1' OR Input1 ='1'  
	ELSE '0' ;             
END ORING;